div_freq_inst : div_freq PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
